package eth_reg_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;


  class class_name extends uvm_reg;
  endclass

  
endpackage
