module top;


  
endmodule
